sin,sina,sitt
henne
hans
